wewerwerwer