Address geneneration unit