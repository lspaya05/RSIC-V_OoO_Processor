//Name: Leonard Paya
//Date: 09/08/2025

// This is the package for the general purpose 32-bit RISC-V processor. It contains the 
//  needed instructions and functions for the following Instruction sets:
//  -   RV32I: Integer
//  -   RV32M: Integer Multiplication and Division
//  -   RV32A: Atomic Instructions
//  -   RV32F: Single Precision Floating Point 
//  -   RV32D: Double Precision Floating Point

// Source: "The RISC-V Instruction Set Manual Volume I: Unprivileged ISA"
// Link: https://riscv.atlassian.net/wiki/spaces/HOME/pages/16154769/RISC-V+Technical+Specifications
// Version: 20250508
// Published: May 2025

package RV32G;
    import RV32I::*;
    import RV32M::*;
    import RV32A::*;
    import RV32F::*;
    import RV32D::*;
endpackage