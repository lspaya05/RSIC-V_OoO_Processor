// Name: Leonard Paya
// Date: 11/20/2025
