//Name: Leonard Paya
//Date: 09/08/2025

//  

// Source: "The RISC-V Instruction Set Manual Volume I: Unprivileged ISA"
// Link: https://riscv.atlassian.net/wiki/spaces/HOME/pages/16154769/RISC-V+Technical+Specifications
// Version: 20250508
// Published: May 2025

package RV32F;

endpackage