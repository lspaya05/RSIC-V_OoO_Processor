// Name: Leonard Paya
// Date: 

module ALU_FP #( 
    parameter 
);

endmodule